`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.11.2018 16:57:00
// Design Name: 
// Module Name: test_bench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module test_bench;

	// Inputs
	reg clk,reset;
	reg [31:0] a;
	reg [31:0] b;

	// Outputs
	wire [31:0] fprod;

	// Instantiate the Unit Under Test (UUT)
	fpmul uut ( 
		.clk(clk), 
		.reset(reset),
		.a(a),
		.b(b),
		.fprod(fprod)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		a = 0;
		b = 0;

		// Wait 100 ns for global reset to finish
		#100;
        	clk = 0;//01000001101010010100011110101110==21.16
		a = 32'b11000000100100110011001100110011;//-4.6;
		b = 32'b11000000100100110011001100110011;//-4.6
		// Add stimulus here
#200;
		    	clk = 0;//11000000001100001010001111010111==-2.76
		a = 32'b11000000100100110011001100110011;//-4.6;
		b = 32'b00111111000110011001100110011010;//0.6
		// Add stimulus here
#300;

    	clk = 0;//10111111111101011100001010001111==-1.92
		a = 32'b01000000010011001100110011001101;//3.2;
		b = 32'b10111111000110011001100110011010;//-0.6
		// Add stimulus here
#400;
 	clk = 0;//01001010100101010000111101101110==4884407.0
		a = 32'b01000101000010100111000011001101;//2215.05;
		b = 32'b01000101000010011101000110011010;//2205.10
		// Add stimulus here
#500;
	end	
     always #50 clk=(~clk);  
endmodule
